module vape

import (
	net.http
)

pub struct Context {
pub:
	request http.Request
}
